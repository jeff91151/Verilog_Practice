module top_module (
    input clk,
    input reset,     // synchronous reset
    input w,
    output z);

    parameter A = 0, B = 1, C = 2, D = 3, E = 4, F = 5;
    reg [2:0] next_state, state;
    
    always @(*) begin
       
        case (state)
            A: next_state = w ? B : A ;
            B: next_state = w ? C : D ;
            C: next_state = w ? E : D ;
            D: next_state = w ? F : A ;
            E: next_state = w ? E : D ;
            F: next_state = w ? C : D ;
        endcase
        
    end
    always @(posedge clk) begin
        
        if (reset) begin
           state <= A; 
        end else begin
           state <= next_state; 
        end
    end
    assign z = (state == E)||(state == F);
    
endmodule
